// Create Date: 12/07/2024 09:01:25 PM
// Design Name: 
// Module Name: timer_count_dw_clk4_test
// Project Name: 
// 
//////////////////////////////////////////////////////////////////////////////////


module timer_count_dw_clk4_test;
    
endmodule